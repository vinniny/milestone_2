`timescale 1ns/1ps
// Immediate generator for RV32I
module immgen (
    input  logic [31:0] instr,
    output logic [31:0] imm_i,
    output logic [31:0] imm_s,
    output logic [31:0] imm_b,
    output logic [31:0] imm_u,
    output logic [31:0] imm_j
);
    // Stub
endmodule

