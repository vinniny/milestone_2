`timescale 1ns/1ps
// Branch comparator
module brc (
    input  logic [31:0] rs1,
    input  logic [31:0] rs2,
    input  logic [2:0]  funct3,   // branch type
    output logic        take      // 1 if branch taken
);
    // Stub
endmodule

