`timescale 1ns/1ps
// Instruction memory interface (simple ROM-like)
module imem (
    input  logic        clk,
    input  logic [31:0] addr,
    output logic [31:0] rdata
);
    // Stub
endmodule

