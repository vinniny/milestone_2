`timescale 1ns/1ps
// Program counter register
module pc (
    input  logic        clk,
    input  logic        rst,
    input  logic [31:0] pc_next,
    output logic [31:0] pc_curr
);
    // Stub
endmodule

